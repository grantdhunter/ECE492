// niosII_system.v

// Generated using ACDS version 12.1sp1 243 at 2014.02.11.10:45:36

`timescale 1 ps / 1 ps
module niosII_system (
		input  wire        clk_0_clk_in_clk,                 //              clk_0_clk_in.clk
		input  wire        clk_0_clk_in_reset_reset_n,       //        clk_0_clk_in_reset.reset_n
		output wire [11:0] sdram_0_wire_addr,                //              sdram_0_wire.addr
		output wire [1:0]  sdram_0_wire_ba,                  //                          .ba
		output wire        sdram_0_wire_cas_n,               //                          .cas_n
		output wire        sdram_0_wire_cke,                 //                          .cke
		output wire        sdram_0_wire_cs_n,                //                          .cs_n
		inout  wire [15:0] sdram_0_wire_dq,                  //                          .dq
		output wire [1:0]  sdram_0_wire_dqm,                 //                          .dqm
		output wire        sdram_0_wire_ras_n,               //                          .ras_n
		output wire        sdram_0_wire_we_n,                //                          .we_n
		input  wire        pio_0_external_connection_export  // pio_0_external_connection.export
	);

	wire         altpll_0_c1_clk;                                                                                     // altpll_0:c1 -> [addr_router:clk, addr_router_001:clk, altpll_0:clk, burst_adapter:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, crosser:in_clk, crosser_001:in_clk, crosser_002:in_clk, crosser_003:out_clk, crosser_004:out_clk, crosser_005:out_clk, id_router:clk, id_router_001:clk, id_router_005:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, leds:clk, leds_s1_translator:clk, leds_s1_translator_avalon_universal_slave_0_agent:clk, leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, nios2_qsys_0:clk, nios2_qsys_0_data_master_translator:clk, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_0_instruction_master_translator:clk, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_0_jtag_debug_module_translator:clk, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_005:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller:clk, sdram_0:clk, sdram_0_s1_translator:clk, sdram_0_s1_translator_avalon_universal_slave_0_agent:clk, sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter:clk, width_adapter_001:clk]
	wire         altpll_0_c0_clk;                                                                                     // altpll_0:c0 -> [crosser:out_clk, crosser_001:out_clk, crosser_002:out_clk, crosser_003:in_clk, crosser_004:in_clk, crosser_005:in_clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, jtag_uart_0:clk, jtag_uart_0_avalon_jtag_slave_translator:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rst_controller_001:clk, sysid_qsys_0:clock, sysid_qsys_0_control_slave_translator:clk, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:clk, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer_0:clk, timer_0_s1_translator:clk, timer_0_s1_translator_avalon_universal_slave_0_agent:clk, timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk]
	wire         nios2_qsys_0_data_master_waitrequest;                                                                // nios2_qsys_0_data_master_translator:av_waitrequest -> nios2_qsys_0:d_waitrequest
	wire  [31:0] nios2_qsys_0_data_master_writedata;                                                                  // nios2_qsys_0:d_writedata -> nios2_qsys_0_data_master_translator:av_writedata
	wire  [24:0] nios2_qsys_0_data_master_address;                                                                    // nios2_qsys_0:d_address -> nios2_qsys_0_data_master_translator:av_address
	wire         nios2_qsys_0_data_master_write;                                                                      // nios2_qsys_0:d_write -> nios2_qsys_0_data_master_translator:av_write
	wire         nios2_qsys_0_data_master_read;                                                                       // nios2_qsys_0:d_read -> nios2_qsys_0_data_master_translator:av_read
	wire  [31:0] nios2_qsys_0_data_master_readdata;                                                                   // nios2_qsys_0_data_master_translator:av_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_debugaccess;                                                                // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_0_data_master_translator:av_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                                                                 // nios2_qsys_0:d_byteenable -> nios2_qsys_0_data_master_translator:av_byteenable
	wire         nios2_qsys_0_instruction_master_waitrequest;                                                         // nios2_qsys_0_instruction_master_translator:av_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [24:0] nios2_qsys_0_instruction_master_address;                                                             // nios2_qsys_0:i_address -> nios2_qsys_0_instruction_master_translator:av_address
	wire         nios2_qsys_0_instruction_master_read;                                                                // nios2_qsys_0:i_read -> nios2_qsys_0_instruction_master_translator:av_read
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                                                            // nios2_qsys_0_instruction_master_translator:av_readdata -> nios2_qsys_0:i_readdata
	wire   [1:0] leds_s1_translator_avalon_anti_slave_0_address;                                                      // leds_s1_translator:av_address -> leds:address
	wire  [31:0] leds_s1_translator_avalon_anti_slave_0_readdata;                                                     // leds:readdata -> leds_s1_translator:av_readdata
	wire         sdram_0_s1_translator_avalon_anti_slave_0_waitrequest;                                               // sdram_0:za_waitrequest -> sdram_0_s1_translator:av_waitrequest
	wire  [15:0] sdram_0_s1_translator_avalon_anti_slave_0_writedata;                                                 // sdram_0_s1_translator:av_writedata -> sdram_0:az_data
	wire  [21:0] sdram_0_s1_translator_avalon_anti_slave_0_address;                                                   // sdram_0_s1_translator:av_address -> sdram_0:az_addr
	wire         sdram_0_s1_translator_avalon_anti_slave_0_chipselect;                                                // sdram_0_s1_translator:av_chipselect -> sdram_0:az_cs
	wire         sdram_0_s1_translator_avalon_anti_slave_0_write;                                                     // sdram_0_s1_translator:av_write -> sdram_0:az_wr_n
	wire         sdram_0_s1_translator_avalon_anti_slave_0_read;                                                      // sdram_0_s1_translator:av_read -> sdram_0:az_rd_n
	wire  [15:0] sdram_0_s1_translator_avalon_anti_slave_0_readdata;                                                  // sdram_0:za_data -> sdram_0_s1_translator:av_readdata
	wire         sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid;                                             // sdram_0:za_valid -> sdram_0_s1_translator:av_readdatavalid
	wire   [1:0] sdram_0_s1_translator_avalon_anti_slave_0_byteenable;                                                // sdram_0_s1_translator:av_byteenable -> sdram_0:az_be_n
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_writedata;                                                 // timer_0_s1_translator:av_writedata -> timer_0:writedata
	wire   [2:0] timer_0_s1_translator_avalon_anti_slave_0_address;                                                   // timer_0_s1_translator:av_address -> timer_0:address
	wire         timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                                // timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	wire         timer_0_s1_translator_avalon_anti_slave_0_write;                                                     // timer_0_s1_translator:av_write -> timer_0:write_n
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_readdata;                                                  // timer_0:readdata -> timer_0_s1_translator:av_readdata
	wire   [0:0] sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address;                                   // sysid_qsys_0_control_slave_translator:av_address -> sysid_qsys_0:address
	wire  [31:0] sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata;                                  // sysid_qsys_0:readdata -> sysid_qsys_0_control_slave_translator:av_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                            // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                              // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire   [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                             // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                  // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                   // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                               // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                             // nios2_qsys_0_jtag_debug_module_translator:av_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire   [8:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                               // nios2_qsys_0_jtag_debug_module_translator:av_address -> nios2_qsys_0:jtag_debug_module_address
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                            // nios2_qsys_0_jtag_debug_module_translator:av_chipselect -> nios2_qsys_0:jtag_debug_module_select
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                 // nios2_qsys_0_jtag_debug_module_translator:av_write -> nios2_qsys_0:jtag_debug_module_write
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                              // nios2_qsys_0:jtag_debug_module_readdata -> nios2_qsys_0_jtag_debug_module_translator:av_readdata
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                         // nios2_qsys_0_jtag_debug_module_translator:av_begintransfer -> nios2_qsys_0:jtag_debug_module_begintransfer
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                           // nios2_qsys_0_jtag_debug_module_translator:av_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                            // nios2_qsys_0_jtag_debug_module_translator:av_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest;                           // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_data_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount;                            // nios2_qsys_0_data_master_translator:uav_burstcount -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata;                             // nios2_qsys_0_data_master_translator:uav_writedata -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [24:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_address;                               // nios2_qsys_0_data_master_translator:uav_address -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock;                                  // nios2_qsys_0_data_master_translator:uav_lock -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_write;                                 // nios2_qsys_0_data_master_translator:uav_write -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_read;                                  // nios2_qsys_0_data_master_translator:uav_read -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata;                              // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_data_master_translator:uav_readdata
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess;                           // nios2_qsys_0_data_master_translator:uav_debugaccess -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable;                            // nios2_qsys_0_data_master_translator:uav_byteenable -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid;                         // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_data_master_translator:uav_readdatavalid
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                    // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_instruction_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount;                     // nios2_qsys_0_instruction_master_translator:uav_burstcount -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata;                      // nios2_qsys_0_instruction_master_translator:uav_writedata -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [24:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address;                        // nios2_qsys_0_instruction_master_translator:uav_address -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock;                           // nios2_qsys_0_instruction_master_translator:uav_lock -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write;                          // nios2_qsys_0_instruction_master_translator:uav_write -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read;                           // nios2_qsys_0_instruction_master_translator:uav_read -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata;                       // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_instruction_master_translator:uav_readdata
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                    // nios2_qsys_0_instruction_master_translator:uav_debugaccess -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable;                     // nios2_qsys_0_instruction_master_translator:uav_byteenable -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                  // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_instruction_master_translator:uav_readdatavalid
	wire         leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // leds_s1_translator:uav_waitrequest -> leds_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // leds_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> leds_s1_translator:uav_burstcount
	wire  [31:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // leds_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> leds_s1_translator:uav_writedata
	wire  [24:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // leds_s1_translator_avalon_universal_slave_0_agent:m0_address -> leds_s1_translator:uav_address
	wire         leds_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // leds_s1_translator_avalon_universal_slave_0_agent:m0_write -> leds_s1_translator:uav_write
	wire         leds_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // leds_s1_translator_avalon_universal_slave_0_agent:m0_lock -> leds_s1_translator:uav_lock
	wire         leds_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // leds_s1_translator_avalon_universal_slave_0_agent:m0_read -> leds_s1_translator:uav_read
	wire  [31:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // leds_s1_translator:uav_readdata -> leds_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // leds_s1_translator:uav_readdatavalid -> leds_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // leds_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> leds_s1_translator:uav_debugaccess
	wire   [3:0] leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // leds_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> leds_s1_translator:uav_byteenable
	wire         leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // leds_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // leds_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // leds_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // leds_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> leds_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // leds_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> leds_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // sdram_0_s1_translator:uav_waitrequest -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [1:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_0_s1_translator:uav_burstcount
	wire  [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_0_s1_translator:uav_writedata
	wire  [24:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_0_s1_translator:uav_address
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_0_s1_translator:uav_write
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_0_s1_translator:uav_lock
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_0_s1_translator:uav_read
	wire  [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // sdram_0_s1_translator:uav_readdata -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // sdram_0_s1_translator:uav_readdatavalid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_0_s1_translator:uav_debugaccess
	wire   [1:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_0_s1_translator:uav_byteenable
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [80:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [80:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [15:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	wire  [24:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	wire   [3:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                           // timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                            // timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // sysid_qsys_0_control_slave_translator:uav_waitrequest -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_qsys_0_control_slave_translator:uav_burstcount
	wire  [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                   // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_qsys_0_control_slave_translator:uav_writedata
	wire  [24:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                     // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_qsys_0_control_slave_translator:uav_address
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_qsys_0_control_slave_translator:uav_write
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                        // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_qsys_0_control_slave_translator:uav_lock
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                        // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_qsys_0_control_slave_translator:uav_read
	wire  [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                    // sysid_qsys_0_control_slave_translator:uav_readdata -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // sysid_qsys_0_control_slave_translator:uav_readdatavalid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_qsys_0_control_slave_translator:uav_debugaccess
	wire   [3:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_qsys_0_control_slave_translator:uav_byteenable
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                 // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;           // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;            // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;           // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire  [24:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // nios2_qsys_0_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_0_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;               // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_0_jtag_debug_module_translator:uav_writedata
	wire  [24:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                 // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_0_jtag_debug_module_translator:uav_address
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_0_jtag_debug_module_translator:uav_write
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_0_jtag_debug_module_translator:uav_lock
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_0_jtag_debug_module_translator:uav_read
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                // nios2_qsys_0_jtag_debug_module_translator:uav_readdata -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // nios2_qsys_0_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_0_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_0_jtag_debug_module_translator:uav_byteenable
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;            // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [98:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;            // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [98:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                  // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                        // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [97:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                         // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                        // addr_router:sink_ready -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;           // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                 // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;         // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [97:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                  // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                 // addr_router_001:sink_ready -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // leds_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         leds_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // leds_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // leds_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [97:0] leds_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // leds_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         leds_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router:sink_ready -> leds_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [79:0] sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_001:sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [97:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_002:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                       // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [97:0] sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                        // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_003:sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [97:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_004:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [97:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_005:sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         burst_adapter_source0_endofpacket;                                                                   // burst_adapter:source0_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         burst_adapter_source0_valid;                                                                         // burst_adapter:source0_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         burst_adapter_source0_startofpacket;                                                                 // burst_adapter:source0_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [79:0] burst_adapter_source0_data;                                                                          // burst_adapter:source0_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire         burst_adapter_source0_ready;                                                                         // sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [5:0] burst_adapter_source0_channel;                                                                       // burst_adapter:source0_channel -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rst_controller_reset_out_reset;                                                                      // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, altpll_0:reset, burst_adapter:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, crosser:in_reset, crosser_001:in_reset, crosser_002:in_reset, crosser_003:out_reset, crosser_004:out_reset, crosser_005:out_reset, id_router:reset, id_router_001:reset, id_router_005:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, leds:reset_n, leds_s1_translator:reset, leds_s1_translator_avalon_universal_slave_0_agent:reset, leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, nios2_qsys_0:reset_n, nios2_qsys_0_data_master_translator:reset, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_instruction_master_translator:reset, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_005:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sdram_0:reset_n, sdram_0_s1_translator:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                                                          // nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                                                  // rst_controller_001:reset_out -> [crosser:out_reset, crosser_001:out_reset, crosser_002:out_reset, crosser_003:in_reset, crosser_004:in_reset, crosser_005:in_reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, sysid_qsys_0:reset_n, sysid_qsys_0_control_slave_translator:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0:reset_n, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         cmd_xbar_demux_src0_endofpacket;                                                                     // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                           // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                   // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src0_data;                                                                            // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [5:0] cmd_xbar_demux_src0_channel;                                                                         // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                           // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                     // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                           // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                   // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [97:0] cmd_xbar_demux_src1_data;                                                                            // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire   [5:0] cmd_xbar_demux_src1_channel;                                                                         // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                           // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                                 // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                       // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                               // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src0_data;                                                                        // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [5:0] cmd_xbar_demux_001_src0_channel;                                                                     // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                       // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                                 // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                       // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                               // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src1_data;                                                                        // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire   [5:0] cmd_xbar_demux_001_src1_channel;                                                                     // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                       // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                                 // cmd_xbar_demux_001:src2_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                       // cmd_xbar_demux_001:src2_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                               // cmd_xbar_demux_001:src2_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_demux_001_src2_data;                                                                        // cmd_xbar_demux_001:src2_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [5:0] cmd_xbar_demux_001_src2_channel;                                                                     // cmd_xbar_demux_001:src2_channel -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                     // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                           // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                   // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [97:0] rsp_xbar_demux_src0_data;                                                                            // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [5:0] rsp_xbar_demux_src0_channel;                                                                         // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                           // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                     // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                           // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                   // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [97:0] rsp_xbar_demux_src1_data;                                                                            // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [5:0] rsp_xbar_demux_src1_channel;                                                                         // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                           // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                                 // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                       // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                               // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [97:0] rsp_xbar_demux_001_src0_data;                                                                        // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [5:0] rsp_xbar_demux_001_src0_channel;                                                                     // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                       // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                                 // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                       // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                               // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [97:0] rsp_xbar_demux_001_src1_data;                                                                        // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire   [5:0] rsp_xbar_demux_001_src1_channel;                                                                     // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                       // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                                 // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                       // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                               // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [97:0] rsp_xbar_demux_005_src0_data;                                                                        // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink2_data
	wire   [5:0] rsp_xbar_demux_005_src0_channel;                                                                     // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                       // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_005:src0_ready
	wire         addr_router_src_endofpacket;                                                                         // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                               // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                                       // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [97:0] addr_router_src_data;                                                                                // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [5:0] addr_router_src_channel;                                                                             // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                               // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                        // rsp_xbar_mux:src_endofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                              // rsp_xbar_mux:src_valid -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                      // rsp_xbar_mux:src_startofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [97:0] rsp_xbar_mux_src_data;                                                                               // rsp_xbar_mux:src_data -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [5:0] rsp_xbar_mux_src_channel;                                                                            // rsp_xbar_mux:src_channel -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_src_ready;                                                                              // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire         addr_router_001_src_endofpacket;                                                                     // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         addr_router_001_src_valid;                                                                           // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire         addr_router_001_src_startofpacket;                                                                   // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [97:0] addr_router_001_src_data;                                                                            // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [5:0] addr_router_001_src_channel;                                                                         // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire         addr_router_001_src_ready;                                                                           // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                    // rsp_xbar_mux_001:src_endofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                          // rsp_xbar_mux_001:src_valid -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                  // rsp_xbar_mux_001:src_startofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [97:0] rsp_xbar_mux_001_src_data;                                                                           // rsp_xbar_mux_001:src_data -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [5:0] rsp_xbar_mux_001_src_channel;                                                                        // rsp_xbar_mux_001:src_channel -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                          // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                        // cmd_xbar_mux:src_endofpacket -> leds_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                              // cmd_xbar_mux:src_valid -> leds_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                      // cmd_xbar_mux:src_startofpacket -> leds_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] cmd_xbar_mux_src_data;                                                                               // cmd_xbar_mux:src_data -> leds_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [5:0] cmd_xbar_mux_src_channel;                                                                            // cmd_xbar_mux:src_channel -> leds_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                              // leds_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                           // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                                 // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                         // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [97:0] id_router_src_data;                                                                                  // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [5:0] id_router_src_channel;                                                                               // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                                 // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         crosser_out_ready;                                                                                   // timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire         id_router_002_src_endofpacket;                                                                       // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                             // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                     // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [97:0] id_router_002_src_data;                                                                              // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [5:0] id_router_002_src_channel;                                                                           // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                             // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         crosser_001_out_ready;                                                                               // sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_001:out_ready
	wire         id_router_003_src_endofpacket;                                                                       // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                             // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                     // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [97:0] id_router_003_src_data;                                                                              // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [5:0] id_router_003_src_channel;                                                                           // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                             // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         crosser_002_out_ready;                                                                               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_002:out_ready
	wire         id_router_004_src_endofpacket;                                                                       // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                             // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                     // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [97:0] id_router_004_src_data;                                                                              // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [5:0] id_router_004_src_channel;                                                                           // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                             // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_001_src2_ready;                                                                       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	wire         id_router_005_src_endofpacket;                                                                       // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                             // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                     // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [97:0] id_router_005_src_data;                                                                              // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [5:0] id_router_005_src_channel;                                                                           // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                             // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                    // cmd_xbar_mux_001:src_endofpacket -> width_adapter:in_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                          // cmd_xbar_mux_001:src_valid -> width_adapter:in_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                  // cmd_xbar_mux_001:src_startofpacket -> width_adapter:in_startofpacket
	wire  [97:0] cmd_xbar_mux_001_src_data;                                                                           // cmd_xbar_mux_001:src_data -> width_adapter:in_data
	wire   [5:0] cmd_xbar_mux_001_src_channel;                                                                        // cmd_xbar_mux_001:src_channel -> width_adapter:in_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                          // width_adapter:in_ready -> cmd_xbar_mux_001:src_ready
	wire         width_adapter_src_endofpacket;                                                                       // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire         width_adapter_src_valid;                                                                             // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire         width_adapter_src_startofpacket;                                                                     // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [79:0] width_adapter_src_data;                                                                              // width_adapter:out_data -> burst_adapter:sink0_data
	wire         width_adapter_src_ready;                                                                             // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire   [5:0] width_adapter_src_channel;                                                                           // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire         id_router_001_src_endofpacket;                                                                       // id_router_001:src_endofpacket -> width_adapter_001:in_endofpacket
	wire         id_router_001_src_valid;                                                                             // id_router_001:src_valid -> width_adapter_001:in_valid
	wire         id_router_001_src_startofpacket;                                                                     // id_router_001:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [79:0] id_router_001_src_data;                                                                              // id_router_001:src_data -> width_adapter_001:in_data
	wire   [5:0] id_router_001_src_channel;                                                                           // id_router_001:src_channel -> width_adapter_001:in_channel
	wire         id_router_001_src_ready;                                                                             // width_adapter_001:in_ready -> id_router_001:src_ready
	wire         width_adapter_001_src_endofpacket;                                                                   // width_adapter_001:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         width_adapter_001_src_valid;                                                                         // width_adapter_001:out_valid -> rsp_xbar_demux_001:sink_valid
	wire         width_adapter_001_src_startofpacket;                                                                 // width_adapter_001:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [97:0] width_adapter_001_src_data;                                                                          // width_adapter_001:out_data -> rsp_xbar_demux_001:sink_data
	wire         width_adapter_001_src_ready;                                                                         // rsp_xbar_demux_001:sink_ready -> width_adapter_001:out_ready
	wire   [5:0] width_adapter_001_src_channel;                                                                       // width_adapter_001:out_channel -> rsp_xbar_demux_001:sink_channel
	wire         crosser_out_endofpacket;                                                                             // crosser:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         crosser_out_valid;                                                                                   // crosser:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         crosser_out_startofpacket;                                                                           // crosser:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] crosser_out_data;                                                                                    // crosser:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [5:0] crosser_out_channel;                                                                                 // crosser:out_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src2_endofpacket;                                                                     // cmd_xbar_demux:src2_endofpacket -> crosser:in_endofpacket
	wire         cmd_xbar_demux_src2_valid;                                                                           // cmd_xbar_demux:src2_valid -> crosser:in_valid
	wire         cmd_xbar_demux_src2_startofpacket;                                                                   // cmd_xbar_demux:src2_startofpacket -> crosser:in_startofpacket
	wire  [97:0] cmd_xbar_demux_src2_data;                                                                            // cmd_xbar_demux:src2_data -> crosser:in_data
	wire   [5:0] cmd_xbar_demux_src2_channel;                                                                         // cmd_xbar_demux:src2_channel -> crosser:in_channel
	wire         cmd_xbar_demux_src2_ready;                                                                           // crosser:in_ready -> cmd_xbar_demux:src2_ready
	wire         crosser_001_out_endofpacket;                                                                         // crosser_001:out_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         crosser_001_out_valid;                                                                               // crosser_001:out_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         crosser_001_out_startofpacket;                                                                       // crosser_001:out_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] crosser_001_out_data;                                                                                // crosser_001:out_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [5:0] crosser_001_out_channel;                                                                             // crosser_001:out_channel -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src3_endofpacket;                                                                     // cmd_xbar_demux:src3_endofpacket -> crosser_001:in_endofpacket
	wire         cmd_xbar_demux_src3_valid;                                                                           // cmd_xbar_demux:src3_valid -> crosser_001:in_valid
	wire         cmd_xbar_demux_src3_startofpacket;                                                                   // cmd_xbar_demux:src3_startofpacket -> crosser_001:in_startofpacket
	wire  [97:0] cmd_xbar_demux_src3_data;                                                                            // cmd_xbar_demux:src3_data -> crosser_001:in_data
	wire   [5:0] cmd_xbar_demux_src3_channel;                                                                         // cmd_xbar_demux:src3_channel -> crosser_001:in_channel
	wire         cmd_xbar_demux_src3_ready;                                                                           // crosser_001:in_ready -> cmd_xbar_demux:src3_ready
	wire         crosser_002_out_endofpacket;                                                                         // crosser_002:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         crosser_002_out_valid;                                                                               // crosser_002:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         crosser_002_out_startofpacket;                                                                       // crosser_002:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [97:0] crosser_002_out_data;                                                                                // crosser_002:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [5:0] crosser_002_out_channel;                                                                             // crosser_002:out_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src4_endofpacket;                                                                     // cmd_xbar_demux:src4_endofpacket -> crosser_002:in_endofpacket
	wire         cmd_xbar_demux_src4_valid;                                                                           // cmd_xbar_demux:src4_valid -> crosser_002:in_valid
	wire         cmd_xbar_demux_src4_startofpacket;                                                                   // cmd_xbar_demux:src4_startofpacket -> crosser_002:in_startofpacket
	wire  [97:0] cmd_xbar_demux_src4_data;                                                                            // cmd_xbar_demux:src4_data -> crosser_002:in_data
	wire   [5:0] cmd_xbar_demux_src4_channel;                                                                         // cmd_xbar_demux:src4_channel -> crosser_002:in_channel
	wire         cmd_xbar_demux_src4_ready;                                                                           // crosser_002:in_ready -> cmd_xbar_demux:src4_ready
	wire         crosser_003_out_endofpacket;                                                                         // crosser_003:out_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire         crosser_003_out_valid;                                                                               // crosser_003:out_valid -> rsp_xbar_mux:sink2_valid
	wire         crosser_003_out_startofpacket;                                                                       // crosser_003:out_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [97:0] crosser_003_out_data;                                                                                // crosser_003:out_data -> rsp_xbar_mux:sink2_data
	wire   [5:0] crosser_003_out_channel;                                                                             // crosser_003:out_channel -> rsp_xbar_mux:sink2_channel
	wire         crosser_003_out_ready;                                                                               // rsp_xbar_mux:sink2_ready -> crosser_003:out_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                                 // rsp_xbar_demux_002:src0_endofpacket -> crosser_003:in_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                       // rsp_xbar_demux_002:src0_valid -> crosser_003:in_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                               // rsp_xbar_demux_002:src0_startofpacket -> crosser_003:in_startofpacket
	wire  [97:0] rsp_xbar_demux_002_src0_data;                                                                        // rsp_xbar_demux_002:src0_data -> crosser_003:in_data
	wire   [5:0] rsp_xbar_demux_002_src0_channel;                                                                     // rsp_xbar_demux_002:src0_channel -> crosser_003:in_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                       // crosser_003:in_ready -> rsp_xbar_demux_002:src0_ready
	wire         crosser_004_out_endofpacket;                                                                         // crosser_004:out_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire         crosser_004_out_valid;                                                                               // crosser_004:out_valid -> rsp_xbar_mux:sink3_valid
	wire         crosser_004_out_startofpacket;                                                                       // crosser_004:out_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [97:0] crosser_004_out_data;                                                                                // crosser_004:out_data -> rsp_xbar_mux:sink3_data
	wire   [5:0] crosser_004_out_channel;                                                                             // crosser_004:out_channel -> rsp_xbar_mux:sink3_channel
	wire         crosser_004_out_ready;                                                                               // rsp_xbar_mux:sink3_ready -> crosser_004:out_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                                 // rsp_xbar_demux_003:src0_endofpacket -> crosser_004:in_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                       // rsp_xbar_demux_003:src0_valid -> crosser_004:in_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                               // rsp_xbar_demux_003:src0_startofpacket -> crosser_004:in_startofpacket
	wire  [97:0] rsp_xbar_demux_003_src0_data;                                                                        // rsp_xbar_demux_003:src0_data -> crosser_004:in_data
	wire   [5:0] rsp_xbar_demux_003_src0_channel;                                                                     // rsp_xbar_demux_003:src0_channel -> crosser_004:in_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                       // crosser_004:in_ready -> rsp_xbar_demux_003:src0_ready
	wire         crosser_005_out_endofpacket;                                                                         // crosser_005:out_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire         crosser_005_out_valid;                                                                               // crosser_005:out_valid -> rsp_xbar_mux:sink4_valid
	wire         crosser_005_out_startofpacket;                                                                       // crosser_005:out_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [97:0] crosser_005_out_data;                                                                                // crosser_005:out_data -> rsp_xbar_mux:sink4_data
	wire   [5:0] crosser_005_out_channel;                                                                             // crosser_005:out_channel -> rsp_xbar_mux:sink4_channel
	wire         crosser_005_out_ready;                                                                               // rsp_xbar_mux:sink4_ready -> crosser_005:out_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                                 // rsp_xbar_demux_004:src0_endofpacket -> crosser_005:in_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                       // rsp_xbar_demux_004:src0_valid -> crosser_005:in_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                               // rsp_xbar_demux_004:src0_startofpacket -> crosser_005:in_startofpacket
	wire  [97:0] rsp_xbar_demux_004_src0_data;                                                                        // rsp_xbar_demux_004:src0_data -> crosser_005:in_data
	wire   [5:0] rsp_xbar_demux_004_src0_channel;                                                                     // rsp_xbar_demux_004:src0_channel -> crosser_005:in_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                       // crosser_005:in_ready -> rsp_xbar_demux_004:src0_ready
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                                                              // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         irq_mapper_receiver0_irq;                                                                            // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                                                       // timer_0:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                                                            // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                                                   // jtag_uart_0:av_irq -> irq_synchronizer_001:receiver_irq

	niosII_system_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (altpll_0_c1_clk),                                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                             //                   reset_n.reset_n
		.d_address                             (nios2_qsys_0_data_master_address),                                            //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                               //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                                              //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                                          //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                                        //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                                 //                          .waitrequest
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                                  //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                             // custom_instruction_master.readra
	);

	niosII_system_leds leds (
		.clk      (altpll_0_c1_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address  (leds_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (leds_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (pio_0_external_connection_export)                 // external_connection.export
	);

	niosII_system_sdram_0 sdram_0 (
		.clk            (altpll_0_c1_clk),                                         //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                         // reset.reset_n
		.az_addr        (sdram_0_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_0_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_0_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_0_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_0_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_0_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_0_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_0_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_0_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_0_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_0_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_0_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_0_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_0_wire_dq),                                         //      .export
		.zs_dqm         (sdram_0_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_0_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_0_wire_we_n)                                        //      .export
	);

	niosII_system_altpll_0 altpll_0 (
		.clk       (altpll_0_c1_clk),                //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset), // inclk_interface_reset.reset
		.read      (),                               //             pll_slave.read
		.write     (),                               //                      .write
		.address   (),                               //                      .address
		.readdata  (),                               //                      .readdata
		.writedata (),                               //                      .writedata
		.c0        (altpll_0_c0_clk),                //                    c0.clk
		.c1        (altpll_0_c1_clk),                //                    c1.clk
		.areset    (),                               //        areset_conduit.export
		.locked    (),                               //        locked_conduit.export
		.phasedone ()                                //     phasedone_conduit.export
	);

	niosII_system_timer_0 timer_0 (
		.clk        (altpll_0_c0_clk),                                      //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                  // reset.reset_n
		.address    (timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)                         //   irq.irq
	);

	niosII_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (altpll_0_c0_clk),                                                    //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                                //         reset.reset_n
		.readdata (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	niosII_system_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_0_c0_clk),                                                          //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                                      //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_001_receiver_irq)                                         //               irq.irq
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) nios2_qsys_0_data_master_translator (
		.clk                   (altpll_0_c1_clk),                                                             //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_qsys_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_qsys_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (nios2_qsys_0_data_master_byteenable),                                         //                          .byteenable
		.av_read               (nios2_qsys_0_data_master_read),                                               //                          .read
		.av_readdata           (nios2_qsys_0_data_master_readdata),                                           //                          .readdata
		.av_write              (nios2_qsys_0_data_master_write),                                              //                          .write
		.av_writedata          (nios2_qsys_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (nios2_qsys_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                        //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                        //               (terminated)
		.av_readdatavalid      (),                                                                            //               (terminated)
		.av_lock               (1'b0),                                                                        //               (terminated)
		.uav_clken             (),                                                                            //               (terminated)
		.av_clken              (1'b1)                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (25),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_0_instruction_master_translator (
		.clk                   (altpll_0_c1_clk),                                                                    //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                     //                     reset.reset
		.uav_address           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_qsys_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_qsys_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (nios2_qsys_0_instruction_master_read),                                               //                          .read
		.av_readdata           (nios2_qsys_0_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount         (1'b1),                                                                               //               (terminated)
		.av_byteenable         (4'b1111),                                                                            //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                                               //               (terminated)
		.av_readdatavalid      (),                                                                                   //               (terminated)
		.av_write              (1'b0),                                                                               //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                               //               (terminated)
		.av_lock               (1'b0),                                                                               //               (terminated)
		.av_debugaccess        (1'b0),                                                                               //               (terminated)
		.uav_clken             (),                                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                                //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) leds_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                    //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (leds_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (leds_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (leds_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (leds_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (leds_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                   //              (terminated)
		.av_read               (),                                                                   //              (terminated)
		.av_writedata          (),                                                                   //              (terminated)
		.av_begintransfer      (),                                                                   //              (terminated)
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_chipselect         (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_0_s1_translator (
		.clk                   (altpll_0_c1_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sdram_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (sdram_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (sdram_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (sdram_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (sdram_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (sdram_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (sdram_0_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (sdram_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_s1_translator (
		.clk                   (altpll_0_c0_clk),                                                       //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                    //                    reset.reset
		.uav_address           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_qsys_0_control_slave_translator (
		.clk                   (altpll_0_c0_clk),                                                                       //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                    //                    reset.reset
		.uav_address           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                                      //              (terminated)
		.av_read               (),                                                                                      //              (terminated)
		.av_writedata          (),                                                                                      //              (terminated)
		.av_begintransfer      (),                                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                                      //              (terminated)
		.av_burstcount         (),                                                                                      //              (terminated)
		.av_byteenable         (),                                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                                      //              (terminated)
		.av_lock               (),                                                                                      //              (terminated)
		.av_chipselect         (),                                                                                      //              (terminated)
		.av_clken              (),                                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                                  //              (terminated)
		.av_debugaccess        (),                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                   (altpll_0_c0_clk),                                                                          //                      clk.clk
		.reset                 (rst_controller_001_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                                         //              (terminated)
		.av_burstcount         (),                                                                                         //              (terminated)
		.av_byteenable         (),                                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                                         //              (terminated)
		.av_lock               (),                                                                                         //              (terminated)
		.av_clken              (),                                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                         //              (terminated)
		.av_outputenable       ()                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (25),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_qsys_0_jtag_debug_module_translator (
		.clk                   (altpll_0_c1_clk),                                                                           //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                                          //              (terminated)
		.av_burstcount         (),                                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                      //              (terminated)
		.av_waitrequest        (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                                          //              (terminated)
		.av_lock               (),                                                                                          //              (terminated)
		.av_clken              (),                                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                                      //              (terminated)
		.av_outputenable       ()                                                                                           //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_BEGIN_BURST           (80),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.PKT_BURST_TYPE_H          (77),
		.PKT_BURST_TYPE_L          (76),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_TRANS_EXCLUSIVE       (66),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_THREAD_ID_H           (88),
		.PKT_THREAD_ID_L           (88),
		.PKT_CACHE_H               (95),
		.PKT_CACHE_L               (92),
		.PKT_DATA_SIDEBAND_H       (79),
		.PKT_DATA_SIDEBAND_L       (79),
		.PKT_QOS_H                 (81),
		.PKT_QOS_L                 (81),
		.PKT_ADDR_SIDEBAND_H       (78),
		.PKT_ADDR_SIDEBAND_L       (78),
		.ST_DATA_W                 (98),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent (
		.clk              (altpll_0_c1_clk),                                                                      //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address       (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_src_valid),                                                               //        rp.valid
		.rp_data          (rsp_xbar_mux_src_data),                                                                //          .data
		.rp_channel       (rsp_xbar_mux_src_channel),                                                             //          .channel
		.rp_startofpacket (rsp_xbar_mux_src_startofpacket),                                                       //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_src_endofpacket),                                                         //          .endofpacket
		.rp_ready         (rsp_xbar_mux_src_ready)                                                                //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_BEGIN_BURST           (80),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.PKT_BURST_TYPE_H          (77),
		.PKT_BURST_TYPE_L          (76),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_TRANS_EXCLUSIVE       (66),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_THREAD_ID_H           (88),
		.PKT_THREAD_ID_L           (88),
		.PKT_CACHE_H               (95),
		.PKT_CACHE_L               (92),
		.PKT_DATA_SIDEBAND_H       (79),
		.PKT_DATA_SIDEBAND_L       (79),
		.PKT_QOS_H                 (81),
		.PKT_QOS_L                 (81),
		.PKT_ADDR_SIDEBAND_H       (78),
		.PKT_ADDR_SIDEBAND_L       (78),
		.ST_DATA_W                 (98),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (4'b0000)
	) nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (altpll_0_c1_clk),                                                                             //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.av_address       (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_001_src_valid),                                                                  //        rp.valid
		.rp_data          (rsp_xbar_mux_001_src_data),                                                                   //          .data
		.rp_channel       (rsp_xbar_mux_001_src_channel),                                                                //          .channel
		.rp_startofpacket (rsp_xbar_mux_001_src_startofpacket),                                                          //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_001_src_endofpacket),                                                            //          .endofpacket
		.rp_ready         (rsp_xbar_mux_001_src_ready)                                                                   //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) leds_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (leds_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (leds_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (leds_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (leds_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (leds_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (leds_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (leds_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (leds_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (leds_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (leds_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (leds_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                     //                .channel
		.rf_sink_ready           (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (leds_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (leds_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (62),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_POSTED          (44),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.PKT_TRANS_LOCK            (47),
		.PKT_SRC_ID_H              (66),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (69),
		.PKT_DEST_ID_L             (67),
		.PKT_BURSTWRAP_H           (54),
		.PKT_BURSTWRAP_L           (52),
		.PKT_BYTE_CNT_H            (51),
		.PKT_BYTE_CNT_L            (49),
		.PKT_PROTECTION_H          (73),
		.PKT_PROTECTION_L          (71),
		.PKT_RESPONSE_STATUS_H     (79),
		.PKT_RESPONSE_STATUS_L     (78),
		.PKT_BURST_SIZE_H          (57),
		.PKT_BURST_SIZE_L          (55),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (80),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sdram_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                     //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                     //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                      //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                               //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                   //                .channel
		.rf_sink_ready           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (81),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                               //              cp.ready
		.cp_valid                (crosser_out_valid),                                                               //                .valid
		.cp_data                 (crosser_out_data),                                                                //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                         //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                             //                .channel
		.rf_sink_ready           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                        // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                     // (terminated)
		.csr_read          (1'b0),                                                                      // (terminated)
		.csr_write         (1'b0),                                                                      // (terminated)
		.csr_readdata      (),                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                      // (terminated)
		.almost_full_data  (),                                                                          // (terminated)
		.almost_empty_data (),                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                      // (terminated)
		.out_startofpacket (),                                                                          // (terminated)
		.out_endofpacket   (),                                                                          // (terminated)
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_channel        (1'b0),                                                                      // (terminated)
		.out_channel       ()                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_001_out_ready),                                                                           //              cp.ready
		.cp_valid                (crosser_001_out_valid),                                                                           //                .valid
		.cp_data                 (crosser_001_out_data),                                                                            //                .data
		.cp_startofpacket        (crosser_001_out_startofpacket),                                                                   //                .startofpacket
		.cp_endofpacket          (crosser_001_out_endofpacket),                                                                     //                .endofpacket
		.cp_channel              (crosser_001_out_channel),                                                                         //                .channel
		.rf_sink_ready           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                                           //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                                      // (terminated)
		.out_startofpacket (),                                                                                          // (terminated)
		.out_endofpacket   (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c0_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_002_out_ready),                                                                              //              cp.ready
		.cp_valid                (crosser_002_out_valid),                                                                              //                .valid
		.cp_data                 (crosser_002_out_data),                                                                               //                .data
		.cp_startofpacket        (crosser_002_out_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (crosser_002_out_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (crosser_002_out_channel),                                                                            //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c0_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (32),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_0_c0_clk),                                                                              //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                                         // (terminated)
		.out_startofpacket (),                                                                                             // (terminated)
		.out_endofpacket   (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (60),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (61),
		.PKT_TRANS_POSTED          (62),
		.PKT_TRANS_WRITE           (63),
		.PKT_TRANS_READ            (64),
		.PKT_TRANS_LOCK            (65),
		.PKT_SRC_ID_H              (84),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (87),
		.PKT_DEST_ID_L             (85),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (67),
		.PKT_PROTECTION_H          (91),
		.PKT_PROTECTION_L          (89),
		.PKT_RESPONSE_STATUS_H     (97),
		.PKT_RESPONSE_STATUS_L     (96),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (98),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_0_c1_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src2_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src2_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_001_src2_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src2_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src2_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src2_channel),                                                                     //                .channel
		.rf_sink_ready           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (99),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_0_c1_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	niosII_system_addr_router addr_router (
		.sink_ready         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_src_valid),                                                                //          .valid
		.src_data           (addr_router_src_data),                                                                 //          .data
		.src_channel        (addr_router_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                           //          .endofpacket
	);

	niosII_system_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                                   //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                                   //          .valid
		.src_data           (addr_router_001_src_data),                                                                    //          .data
		.src_channel        (addr_router_001_src_channel),                                                                 //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                              //          .endofpacket
	);

	niosII_system_id_router id_router (
		.sink_ready         (leds_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (leds_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (leds_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (leds_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (leds_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                //       src.ready
		.src_valid          (id_router_src_valid),                                                //          .valid
		.src_data           (id_router_src_data),                                                 //          .data
		.src_channel        (id_router_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                           //          .endofpacket
	);

	niosII_system_id_router_001 id_router_001 (
		.sink_ready         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                               //       src.ready
		.src_valid          (id_router_001_src_valid),                                               //          .valid
		.src_data           (id_router_001_src_data),                                                //          .data
		.src_channel        (id_router_001_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                          //          .endofpacket
	);

	niosII_system_id_router_002 id_router_002 (
		.sink_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                               //       src.ready
		.src_valid          (id_router_002_src_valid),                                               //          .valid
		.src_data           (id_router_002_src_data),                                                //          .data
		.src_channel        (id_router_002_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                          //          .endofpacket
	);

	niosII_system_id_router_002 id_router_003 (
		.sink_ready         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                               //       src.ready
		.src_valid          (id_router_003_src_valid),                                                               //          .valid
		.src_data           (id_router_003_src_data),                                                                //          .data
		.src_channel        (id_router_003_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                          //          .endofpacket
	);

	niosII_system_id_router_002 id_router_004 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c0_clk),                                                                          //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_004_src_valid),                                                                  //          .valid
		.src_data           (id_router_004_src_data),                                                                   //          .data
		.src_channel        (id_router_004_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                             //          .endofpacket
	);

	niosII_system_id_router_005 id_router_005 (
		.sink_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_0_c1_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                   //          .valid
		.src_data           (id_router_005_src_data),                                                                    //          .data
		.src_channel        (id_router_005_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                              //          .endofpacket
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (42),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (62),
		.PKT_BYTE_CNT_H            (51),
		.PKT_BYTE_CNT_L            (49),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (57),
		.PKT_BURST_SIZE_L          (55),
		.PKT_BURST_TYPE_H          (59),
		.PKT_BURST_TYPE_L          (58),
		.PKT_BURSTWRAP_H           (54),
		.PKT_BURSTWRAP_L           (52),
		.PKT_TRANS_COMPRESSED_READ (43),
		.PKT_TRANS_WRITE           (45),
		.PKT_TRANS_READ            (46),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (80),
		.ST_CHANNEL_W              (6),
		.OUT_BYTE_CNT_H            (50),
		.OUT_BURSTWRAP_H           (54),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (altpll_0_c1_clk),                     //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~clk_0_clk_in_reset_reset_n),                // reset_in0.reset
		.reset_in1  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (altpll_0_c1_clk),                            //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~clk_0_clk_in_reset_reset_n),                // reset_in0.reset
		.reset_in1  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (altpll_0_c0_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),         // reset_out.reset
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	niosII_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (altpll_0_c1_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket),   //          .endofpacket
		.src4_ready         (cmd_xbar_demux_src4_ready),         //      src4.ready
		.src4_valid         (cmd_xbar_demux_src4_valid),         //          .valid
		.src4_data          (cmd_xbar_demux_src4_data),          //          .data
		.src4_channel       (cmd_xbar_demux_src4_channel),       //          .channel
		.src4_startofpacket (cmd_xbar_demux_src4_startofpacket), //          .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_src4_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_001_src_ready),             //      sink.ready
		.sink_channel       (addr_router_001_src_channel),           //          .channel
		.sink_data          (addr_router_001_src_data),              //          .data
		.sink_startofpacket (addr_router_001_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_001_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_001_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (altpll_0_c1_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (altpll_0_c1_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (altpll_0_c1_clk),                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),         //          .channel
		.sink_data          (width_adapter_001_src_data),            //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (altpll_0_c0_clk),                       //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_demux_002 rsp_xbar_demux_005 (
		.clk                (altpll_0_c1_clk),                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	niosII_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (altpll_0_c1_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (crosser_003_out_ready),                 //     sink2.ready
		.sink2_valid         (crosser_003_out_valid),                 //          .valid
		.sink2_channel       (crosser_003_out_channel),               //          .channel
		.sink2_data          (crosser_003_out_data),                  //          .data
		.sink2_startofpacket (crosser_003_out_startofpacket),         //          .startofpacket
		.sink2_endofpacket   (crosser_003_out_endofpacket),           //          .endofpacket
		.sink3_ready         (crosser_004_out_ready),                 //     sink3.ready
		.sink3_valid         (crosser_004_out_valid),                 //          .valid
		.sink3_channel       (crosser_004_out_channel),               //          .channel
		.sink3_data          (crosser_004_out_data),                  //          .data
		.sink3_startofpacket (crosser_004_out_startofpacket),         //          .startofpacket
		.sink3_endofpacket   (crosser_004_out_endofpacket),           //          .endofpacket
		.sink4_ready         (crosser_005_out_ready),                 //     sink4.ready
		.sink4_valid         (crosser_005_out_valid),                 //          .valid
		.sink4_channel       (crosser_005_out_channel),               //          .channel
		.sink4_data          (crosser_005_out_data),                  //          .data
		.sink4_startofpacket (crosser_005_out_startofpacket),         //          .startofpacket
		.sink4_endofpacket   (crosser_005_out_endofpacket)            //          .endofpacket
	);

	niosII_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (altpll_0_c1_clk),                       //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_005_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (60),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (69),
		.IN_PKT_BYTE_CNT_L             (67),
		.IN_PKT_TRANS_COMPRESSED_READ  (61),
		.IN_PKT_BURSTWRAP_H            (72),
		.IN_PKT_BURSTWRAP_L            (70),
		.IN_PKT_BURST_SIZE_H           (75),
		.IN_PKT_BURST_SIZE_L           (73),
		.IN_PKT_RESPONSE_STATUS_H      (97),
		.IN_PKT_RESPONSE_STATUS_L      (96),
		.IN_PKT_TRANS_EXCLUSIVE        (66),
		.IN_PKT_BURST_TYPE_H           (77),
		.IN_PKT_BURST_TYPE_L           (76),
		.IN_ST_DATA_W                  (98),
		.OUT_PKT_ADDR_H                (42),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (51),
		.OUT_PKT_BYTE_CNT_L            (49),
		.OUT_PKT_TRANS_COMPRESSED_READ (43),
		.OUT_PKT_BURST_SIZE_H          (57),
		.OUT_PKT_BURST_SIZE_L          (55),
		.OUT_PKT_RESPONSE_STATUS_H     (79),
		.OUT_PKT_RESPONSE_STATUS_L     (78),
		.OUT_PKT_TRANS_EXCLUSIVE       (48),
		.OUT_PKT_BURST_TYPE_H          (59),
		.OUT_PKT_BURST_TYPE_L          (58),
		.OUT_ST_DATA_W                 (80),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (altpll_0_c1_clk),                    //       clk.clk
		.reset                (rst_controller_reset_out_reset),     // clk_reset.reset
		.in_valid             (cmd_xbar_mux_001_src_valid),         //      sink.valid
		.in_channel           (cmd_xbar_mux_001_src_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_mux_001_src_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_mux_001_src_ready),         //          .ready
		.in_data              (cmd_xbar_mux_001_src_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (42),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (51),
		.IN_PKT_BYTE_CNT_L             (49),
		.IN_PKT_TRANS_COMPRESSED_READ  (43),
		.IN_PKT_BURSTWRAP_H            (54),
		.IN_PKT_BURSTWRAP_L            (52),
		.IN_PKT_BURST_SIZE_H           (57),
		.IN_PKT_BURST_SIZE_L           (55),
		.IN_PKT_RESPONSE_STATUS_H      (79),
		.IN_PKT_RESPONSE_STATUS_L      (78),
		.IN_PKT_TRANS_EXCLUSIVE        (48),
		.IN_PKT_BURST_TYPE_H           (59),
		.IN_PKT_BURST_TYPE_L           (58),
		.IN_ST_DATA_W                  (80),
		.OUT_PKT_ADDR_H                (60),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (69),
		.OUT_PKT_BYTE_CNT_L            (67),
		.OUT_PKT_TRANS_COMPRESSED_READ (61),
		.OUT_PKT_BURST_SIZE_H          (75),
		.OUT_PKT_BURST_SIZE_L          (73),
		.OUT_PKT_RESPONSE_STATUS_H     (97),
		.OUT_PKT_RESPONSE_STATUS_L     (96),
		.OUT_PKT_TRANS_EXCLUSIVE       (66),
		.OUT_PKT_BURST_TYPE_H          (77),
		.OUT_PKT_BURST_TYPE_L          (76),
		.OUT_ST_DATA_W                 (98),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (1)
	) width_adapter_001 (
		.clk                  (altpll_0_c1_clk),                     //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_001_src_valid),             //      sink.valid
		.in_channel           (id_router_001_src_channel),           //          .channel
		.in_startofpacket     (id_router_001_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_001_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_001_src_ready),             //          .ready
		.in_data              (id_router_001_src_data),              //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (98),
		.BITS_PER_SYMBOL     (98),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (altpll_0_c1_clk),                    //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),     //  in_clk_reset.reset
		.out_clk           (altpll_0_c0_clk),                    //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset), // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src2_ready),          //            in.ready
		.in_valid          (cmd_xbar_demux_src2_valid),          //              .valid
		.in_startofpacket  (cmd_xbar_demux_src2_startofpacket),  //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src2_endofpacket),    //              .endofpacket
		.in_channel        (cmd_xbar_demux_src2_channel),        //              .channel
		.in_data           (cmd_xbar_demux_src2_data),           //              .data
		.out_ready         (crosser_out_ready),                  //           out.ready
		.out_valid         (crosser_out_valid),                  //              .valid
		.out_startofpacket (crosser_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_out_channel),                //              .channel
		.out_data          (crosser_out_data),                   //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (98),
		.BITS_PER_SYMBOL     (98),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (altpll_0_c1_clk),                    //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),     //  in_clk_reset.reset
		.out_clk           (altpll_0_c0_clk),                    //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset), // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src3_ready),          //            in.ready
		.in_valid          (cmd_xbar_demux_src3_valid),          //              .valid
		.in_startofpacket  (cmd_xbar_demux_src3_startofpacket),  //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src3_endofpacket),    //              .endofpacket
		.in_channel        (cmd_xbar_demux_src3_channel),        //              .channel
		.in_data           (cmd_xbar_demux_src3_data),           //              .data
		.out_ready         (crosser_001_out_ready),              //           out.ready
		.out_valid         (crosser_001_out_valid),              //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),      //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),        //              .endofpacket
		.out_channel       (crosser_001_out_channel),            //              .channel
		.out_data          (crosser_001_out_data),               //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (98),
		.BITS_PER_SYMBOL     (98),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (altpll_0_c1_clk),                    //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),     //  in_clk_reset.reset
		.out_clk           (altpll_0_c0_clk),                    //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset), // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src4_ready),          //            in.ready
		.in_valid          (cmd_xbar_demux_src4_valid),          //              .valid
		.in_startofpacket  (cmd_xbar_demux_src4_startofpacket),  //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src4_endofpacket),    //              .endofpacket
		.in_channel        (cmd_xbar_demux_src4_channel),        //              .channel
		.in_data           (cmd_xbar_demux_src4_data),           //              .data
		.out_ready         (crosser_002_out_ready),              //           out.ready
		.out_valid         (crosser_002_out_valid),              //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),      //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),        //              .endofpacket
		.out_channel       (crosser_002_out_channel),            //              .channel
		.out_data          (crosser_002_out_data),               //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (98),
		.BITS_PER_SYMBOL     (98),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (altpll_0_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c1_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_002_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_002_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_002_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_002_src0_data),          //              .data
		.out_ready         (crosser_003_out_ready),                 //           out.ready
		.out_valid         (crosser_003_out_valid),                 //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_003_out_channel),               //              .channel
		.out_data          (crosser_003_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (98),
		.BITS_PER_SYMBOL     (98),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_004 (
		.in_clk            (altpll_0_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c1_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_003_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_003_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_003_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_003_src0_data),          //              .data
		.out_ready         (crosser_004_out_ready),                 //           out.ready
		.out_valid         (crosser_004_out_valid),                 //              .valid
		.out_startofpacket (crosser_004_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_004_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_004_out_channel),               //              .channel
		.out_data          (crosser_004_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (98),
		.BITS_PER_SYMBOL     (98),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_005 (
		.in_clk            (altpll_0_c0_clk),                       //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_0_c1_clk),                       //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_004_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_004_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_004_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_004_src0_data),          //              .data
		.out_ready         (crosser_005_out_ready),                 //           out.ready
		.out_valid         (crosser_005_out_valid),                 //              .valid
		.out_startofpacket (crosser_005_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_005_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_005_out_channel),               //              .channel
		.out_data          (crosser_005_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	niosII_system_irq_mapper irq_mapper (
		.clk           (altpll_0_c1_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_0_c0_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c1_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (altpll_0_c0_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c1_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

endmodule
