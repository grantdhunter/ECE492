-- German R. Gomez Urbina
-- grgomez@ualberta.ca 

library IEEE;

-- Commonly imported packages:
use IEEE.STD_LOGIC_1164.ALL;
use	IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity adc_tuto is
	port (
		-- 50MHz clock & reset
		CLOCK_50 : in std_logic;
		KEY      : in std_logic_vector(1 downto 0);
		
		-- ADC component
		ADC_SCLK : out std_logic;
		ADC_CS_N : out std_logic;
		ADC_DOUT : in  std_logic;
		ADC_DIN  : out std_logic;
		
		-- SDRAM component
		DRAM_ADDR  : out std_logic_vector(11 downto 0);
		DRAM_BA    : out std_logic_vector(1 downto 0);
		DRAM_CAS_N : out std_logic;
		DRAM_CKE   : out std_logic;
		DRAM_CS_N  : out std_logic;
		DRAM_DQ    : inout std_logic_vector(15 downto 0);
		DRAM_DQM   : out std_logic_vector(1 downto 0);
		DRAM_RAS_N : out std_logic;
		DRAM_WE_N  : out std_logic;
		DRAM_CLK   : out std_logic
		
	);
end adc_tuto;

architecture structure of adc_tuto is
	 component niosII is
        port (
            clk_clk                                : in    std_logic                     := 'X';             -- clk
            reset_reset_n                          : in    std_logic                     := 'X';             -- reset_n
            de0_nano_adc_0_external_interface_sclk : out   std_logic;                                        -- sclk
            de0_nano_adc_0_external_interface_cs_n : out   std_logic;                                        -- cs_n
            de0_nano_adc_0_external_interface_dout : in    std_logic                     := 'X';             -- dout
            de0_nano_adc_0_external_interface_din  : out   std_logic;                                        -- din
            sdram_0_wire_addr                      : out   std_logic_vector(11 downto 0);                    -- addr
            sdram_0_wire_ba                        : out   std_logic_vector(1 downto 0);                     -- ba
            sdram_0_wire_cas_n                     : out   std_logic;                                        -- cas_n
            sdram_0_wire_cke                       : out   std_logic;                                        -- cke
            sdram_0_wire_cs_n                      : out   std_logic;                                        -- cs_n
            sdram_0_wire_dq                        : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
            sdram_0_wire_dqm                       : out   std_logic_vector(1 downto 0);                     -- dqm
            sdram_0_wire_ras_n                     : out   std_logic;                                        -- ras_n
            sdram_0_wire_we_n                      : out   std_logic;                                        -- we_n
            altpll_0_c0_clk                        : out   std_logic                                         -- clk
        );
    end component niosII;
	
	begin
	u0 : component niosII
        port map (
            clk_clk                                => CLOCK_50,
            reset_reset_n                          => KEY(0),
            de0_nano_adc_0_external_interface_sclk => ADC_SCLK,
            de0_nano_adc_0_external_interface_cs_n => ADC_CS_N,
            de0_nano_adc_0_external_interface_dout => ADC_DOUT,
            de0_nano_adc_0_external_interface_din  => ADC_DIN,
            sdram_0_wire_addr                      => DRAM_ADDR,
            sdram_0_wire_ba                        => DRAM_BA,
            sdram_0_wire_cas_n                     => DRAM_CAS_N,
            sdram_0_wire_cke                       => DRAM_CKE,
            sdram_0_wire_cs_n                      => DRAM_CS_N,
            sdram_0_wire_dq                        => DRAM_DQ,
            sdram_0_wire_dqm                       => DRAM_DQM,
            sdram_0_wire_ras_n                     => DRAM_RAS_N,
            sdram_0_wire_we_n                      => DRAM_WE_N,
            altpll_0_c0_clk                        => DRAM_CLK
        );
end structure;
	
